
module osd_him
  (input clk, rst,
   glip_channel.slave glip_in,
   glip_channel.master glip_out,

   dii_channel.master dii_out,
   dii_channel.slave dii_in);


endmodule // osd_him

