
module osd_scm
  #(parameter VENDORID='x,
    parameter SYSTEMID='x,
    parameter NUM_MOD='x)
   (input clk, rst,
    dii_channel debug_in,
    dii_channel debug_out);
   
   

endmodule
